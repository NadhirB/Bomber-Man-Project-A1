// System-Verilog 'written by Alex Grinshpun May 2018
// New bitmap dudy February 2025
// (c) Technion IIT, Department of Electrical Engineering 2025 



module	playerBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
				   output   logic	[3:0] HitEdgeCode 
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^6 = 64 



 logic	[10:0] HitCodeX ;// offset of Hitcode 
 logic	[10:0] HitCodeY ; 
assign HitCodeX = offsetX >> ( OBJECT_NUMBER_OF_X_BITS - 4 );	// hitedge code MSB of the offset
assign HitCodeY = offsetY >> ( OBJECT_NUMBER_OF_Y_BITS - 4 );	 	 

// generating a smiley bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00;// RGB value in the bitmap representing a transparent pixel 

logic [0:31] [0:31] [7:0] object_colors = {
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h04,8'h04,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h30,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h30,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h0c,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h0c,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00},
	{8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00},
	{8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00},
	{8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h0c,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h0c,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h30,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h30,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h34,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h04,8'h04,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};


//////////--------------------------------------------------------------------------------------------------------------=
//hit bit map has one encoding per edge:  hit_colors[2:0] =   
 
logic [0:15] [0:15] [2:0] hit_colors = 
		  {48'o3333333333333333,     
			48'o1333333333333332,    
			48'o1133333333333322, 
			48'o1113333333333222,
			48'o1111333333332222,
			48'o1111133333322222,
			48'o1111113333222222,
			48'o1111111332222222,
			48'o1111111002222222,
			48'o1111110000222222,
			48'o1111100000022222,
			48'o1111000000002222,
			48'o1110000000000222,
			48'o1100000000000022,
			48'o1000000000000002,
			48'o0000000000000000};

//logic [0:3] [0:3] [3:0] hit_colors = 
//			{16'hc446,
//			 16'h8c62,
//			 16'h8932,
//			 16'h9113};
 
 
// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		HitEdgeCode <= 3'h0;

	end

	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default  
		HitEdgeCode <= 3'h0;

		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket 
			RGBout <= object_colors[offsetY][offsetX];
			HitEdgeCode <= hit_colors[HitCodeY][HitCodeX];	//get hitting edge code from the colors table  
		
		end  	
	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule