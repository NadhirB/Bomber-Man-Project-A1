
// This module is used to generate a letter sequence (a sentence in the same Y coordinates)
// Using a conversion table and 16 letters as parameters we can efficiently use fewer modules to generate more letters

module	letter_sequence	(	
					input	logic	clk,
					input	logic	resetN,
					
					output [4:0] letters [15:0]
 ) ;

 
parameter int num_of_letters = 16;
parameter logic [4:0] letter_0 = 5'd0;
parameter logic [4:0] letter_1 = 5'd0;
parameter logic [4:0] letter_2 = 5'd0;
parameter logic [4:0] letter_3 = 5'd0;
parameter logic [4:0] letter_4 = 5'd0;
parameter logic [4:0] letter_5 = 5'd0;
parameter logic [4:0] letter_6 = 5'd0;
parameter logic [4:0] letter_7 = 5'd0;
parameter logic [4:0] letter_8 = 5'd0;
parameter logic [4:0] letter_9 = 5'd0;
parameter logic [4:0] letter_10 = 5'd0;
parameter logic [4:0] letter_11 = 5'd0;
parameter logic [4:0] letter_12 = 5'd0;
parameter logic [4:0] letter_13 = 5'd0;
parameter logic [4:0] letter_14 = 5'd0;
parameter logic [4:0] letter_15 = 5'd0;



logic [4:0] letters_out [0: num_of_letters - 1];

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		letters_out <= '{5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0 , 5'd0};
	end

	else begin
		letters_out <= '{letter_0, letter_1, letter_2, letter_3, letter_4, letter_5, letter_6, letter_7, letter_8, letter_9, letter_10, letter_11, letter_12, letter_13, letter_14, letter_15};
	end
		
end

assign letters = letters_out ; 

endmodule