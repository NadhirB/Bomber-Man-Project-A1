// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Feb 2025 
//(c) Technion IIT, Department of Electrical Engineering 2025 



module	blastMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket
					input logic [2:0] blast_num,
					input logic blast,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 


localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^5 = 32  everu object 
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 

localparam  int MAZE_NUMBER_OF__X_BITS = 4;  // 2^4 = 16 / /the maze of the objects 
localparam  int MAZE_NUMBER_OF__Y_BITS = 3;  // 2^3 = 8 

//-----

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;
localparam  int MAZE_WIDTH_X = 1 << MAZE_NUMBER_OF__X_BITS ;
localparam  int MAZE_HEIGHT_Y = 1 << MAZE_NUMBER_OF__Y_BITS ;


 logic [10:0] offsetX_LSB  ;
 logic [10:0] offsetY_LSB  ; 
 logic [10:0] offsetX_MSB ;
 logic [10:0] offsetY_MSB  ;
 logic [2:0] blast_num_D;

 assign offsetX_LSB  = offsetX[(TILE_NUMBER_OF_X_BITS-1):0] ; // get lower bits 
 assign offsetY_LSB  = offsetY[(TILE_NUMBER_OF_Y_BITS-1):0] ; // get lower bits 
 assign offsetX_MSB  = offsetX[(TILE_NUMBER_OF_X_BITS + MAZE_NUMBER_OF__X_BITS -1 ):TILE_NUMBER_OF_X_BITS] ; // get higher bits 
 assign offsetY_MSB  = offsetY[(TILE_NUMBER_OF_Y_BITS + MAZE_NUMBER_OF__Y_BITS -1 ):TILE_NUMBER_OF_Y_BITS] ; // get higher bits 
 

 
// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 8 *16 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the understanding 



// This is a Test:

logic [1:0] MazeBitMapMask [0:2] [0:4] [0:4];

logic [1:0] MazeDefaultBitMapMask [0:2] [0:4] [0:4] = '{
	'{'{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b1, 1'b1, 1'b1, 1'b0},			// Regular blast
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0}},
	  
	'{'{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},			// Vertical blast
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0}},
	  
	'{'{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b1, 1'b1, 1'b1, 1'b0},			// Horizontal blast
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0}}};
 

logic [0:TILE_HEIGHT_Y-1] [0:TILE_WIDTH_X-1] [7:0] object_colors = {
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hac,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc4,8'hFF,8'hFF,8'h84,8'hFF,8'h64,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'he4,8'ha0,8'hFF,8'h64,8'hFF,8'h84,8'hFF,8'he4,8'hFF,8'hFF,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'hFF,8'hFF,8'hFF,8'he4,8'hf4,8'he4,8'he4,8'hac,8'hac,8'h64,8'h64,8'he4,8'hf4,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h20,8'hac,8'h64,8'hac,8'hFF,8'hFF,8'hf4,8'hf8,8'hf4,8'hf4,8'h64,8'he4,8'he4,8'hf4,8'hfd,8'h64,8'hFF,8'hFF,8'hac,8'h64,8'hac,8'h8c,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hac,8'h64,8'h84,8'h64,8'h64,8'hac,8'hfe,8'hf8,8'hf0,8'he4,8'he4,8'he4,8'hf4,8'hfd,8'hac,8'h64,8'h64,8'h64,8'h64,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hac,8'h8c,8'hac,8'h64,8'he4,8'hf0,8'hfd,8'hf4,8'hfd,8'hf4,8'he4,8'hfc,8'hfd,8'hf0,8'he4,8'he4,8'h64,8'h64,8'hac,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'h64,8'hac,8'hac,8'he4,8'he4,8'hf4,8'hfd,8'hfd,8'hf4,8'hfd,8'hf0,8'hf4,8'he4,8'hac,8'h64,8'hac,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hf4,8'he4,8'hec,8'h64,8'h84,8'h64,8'he4,8'h84,8'h64,8'he4,8'hf4,8'hfd,8'hfd,8'hfd,8'hfe,8'he4,8'hfc,8'hf4,8'h64,8'hac,8'he4,8'he4,8'h64,8'hFF,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hf4,8'he4,8'hf4,8'ha4,8'hf4,8'h64,8'h64,8'hfd,8'he4,8'hf8,8'hf0,8'hf8,8'hec,8'hf4,8'hfd,8'h64,8'he4,8'he4,8'hf0,8'hf4,8'hfd,8'hec,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'hf4,8'hf4,8'hfe,8'hfe,8'hf4,8'hf4,8'hfd,8'hf4,8'he4,8'hec,8'hf4,8'hec,8'hfc,8'hfd,8'hf8,8'hfd,8'he4,8'h64,8'hfe,8'hfe,8'hf8,8'ha4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'h64,8'h64,8'h64,8'he4,8'hf4,8'hfd,8'hf4,8'hf4,8'hf4,8'hfe,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'he4,8'he4,8'hfd,8'hf8,8'hf0,8'hfc,8'he4,8'he4,8'hFF,8'h84,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h84,8'h64,8'he4,8'hec,8'hfc,8'he4,8'hf4,8'hfc,8'hf4,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'hf8,8'hfe,8'hfe,8'hfe,8'he4,8'he4,8'h64,8'h84,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'h64,8'hac,8'h64,8'h64,8'h64,8'he4,8'he4,8'hf0,8'hf4,8'hfe,8'hfc,8'hf0,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hf0,8'hec,8'hfc,8'hfe,8'hfc,8'he4,8'h84,8'he4,8'h64,8'h64,8'hac,8'hac,8'hFF},
	{8'hFF,8'h8c,8'hac,8'h64,8'h64,8'he4,8'h84,8'he4,8'hf0,8'hfe,8'hfc,8'hec,8'hf4,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hf4,8'hfd,8'hfe,8'hf4,8'hf0,8'he4,8'he4,8'h64,8'h64,8'h64,8'hac,8'h8c,8'hFF},
	{8'hFF,8'hFF,8'h20,8'hFF,8'h64,8'h64,8'he4,8'he4,8'hfe,8'hfd,8'hfe,8'hf4,8'hf4,8'hfd,8'hfd,8'hfe,8'hfc,8'hfd,8'hfc,8'hfd,8'hf4,8'he4,8'hfc,8'he4,8'he4,8'h84,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'h64,8'hFF,8'he4,8'he4,8'hf8,8'hf4,8'hf8,8'hfe,8'he4,8'he4,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfd,8'hf4,8'hf8,8'hf8,8'hfc,8'hf4,8'hec,8'h84,8'h64,8'h64,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'ha4,8'hf8,8'hfd,8'hfe,8'h64,8'he4,8'hfd,8'hf8,8'hfe,8'hfc,8'hec,8'hf0,8'he4,8'he4,8'hf4,8'hfe,8'hf4,8'hf4,8'hfe,8'hfe,8'hf4,8'hf4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'hfd,8'hf4,8'hac,8'he4,8'he4,8'h64,8'hfd,8'hf4,8'hec,8'hf8,8'hf0,8'hf4,8'he4,8'hfd,8'h64,8'h64,8'hf4,8'he4,8'hf4,8'he4,8'hf4,8'hc4,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'ha4,8'he4,8'hFF,8'h64,8'he4,8'he4,8'hac,8'h64,8'hf4,8'hf8,8'he4,8'hfd,8'hfd,8'hfe,8'hfe,8'hf4,8'he4,8'h64,8'hc4,8'he4,8'h64,8'h64,8'h64,8'he4,8'he4,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'h84,8'h64,8'hcc,8'he4,8'hf4,8'hf0,8'hfd,8'hf4,8'hfd,8'hfe,8'hf4,8'he4,8'he4,8'hac,8'h8c,8'h64,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'ha4,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hac,8'hac,8'h84,8'h64,8'he4,8'he4,8'hf0,8'hfd,8'hfc,8'he4,8'hf4,8'hfe,8'hf8,8'hfd,8'hf4,8'he4,8'h84,8'h64,8'h64,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h84,8'h64,8'hac,8'h64,8'h64,8'h8c,8'hfd,8'hf4,8'he4,8'hec,8'he4,8'he4,8'hf8,8'hfe,8'he4,8'h64,8'h64,8'h64,8'h64,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h20,8'hac,8'hac,8'hac,8'hFF,8'hFF,8'h64,8'hfd,8'hf4,8'he4,8'he4,8'h64,8'hf4,8'hf4,8'hf8,8'hf4,8'hFF,8'hFF,8'hac,8'h84,8'h84,8'h8c,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'hFF,8'hFF,8'hFF,8'hFF,8'h84,8'hf4,8'he4,8'h64,8'h64,8'hac,8'h84,8'he4,8'he4,8'hf8,8'hc4,8'hFF,8'hFF,8'hFF,8'h8c,8'h20,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'hFF,8'hFF,8'he4,8'hFF,8'h84,8'hFF,8'h64,8'hFF,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'h84,8'hFF,8'h64,8'hFF,8'hFF,8'ha4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hac,8'hac,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h64,8'h84,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h60,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}};

 
//
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
		blast_num_D <= 0;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		
		if (!blast)
			blast_num_D <= blast_num;		// Charges the last input from the random module
			
		if (InsideRectangle == 1'b1 )	
			begin 
		   	case (MazeBitMapMask[blast_num_D][offsetY_MSB][offsetX_MSB])
					 1'b0 : RGBout <= TRANSPARENT_ENCODING ;
					 1'b1 : RGBout <= object_colors[offsetY_LSB][offsetX_LSB];  
				default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
			end 

	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

