// System-Verilog 'written by Alex Grinshpun May 2018
// New bitmap dudy February 2025
// (c) Technion IIT, Department of Electrical Engineering 2025 



module	playerBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic left_key,
					input logic right_key,
					input logic up_key,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
				   output   logic	[3:0] HitEdgeCode 
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^6 = 64 



 logic	[10:0] HitCodeX ;// offset of Hitcode 
 logic	[10:0] HitCodeY ; 
//assign HitCodeX = offsetX >> ( OBJECT_NUMBER_OF_X_BITS - 2 );	// hitedge code MSB of the offset was 4 and not 2
//assign HitCodeY = offsetY >> ( OBJECT_NUMBER_OF_Y_BITS - 2 );	 	 

// generating a smiley bitmap

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hff;// RGB value in the bitmap representing a transparent pixel 

logic [0:2] [0:31] [0:31] [7:0] object_colors = {
	{{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h46,8'h46,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h46,8'h46,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h46,8'h46,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h46,8'h46,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h65,8'had,8'had,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'had,8'had,8'h65,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'h65,8'had,8'had,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'had,8'had,8'h65,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h46,8'h46,8'hfa,8'hfa,8'hfa,8'hfa,8'h46,8'h46,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h46,8'h46,8'hfa,8'hfa,8'hfa,8'hfa,8'h46,8'h46,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hc5,8'hc5,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hc5,8'hc5,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hfa,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'hfa,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hfa,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'hfa,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}},
	
	{{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff},
	{8'hff,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'hff},
	{8'hff,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'hff},
	{8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff},
	{8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}},
	
	{{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65},
	{8'hff,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65},
	{8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h65,8'h65,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'h65,8'h65,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'h65,8'h65,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'h65,8'h65,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff}}
	
	};


//////////--------------------------------------------------------------------------------------------------------------=
//hit bit map has one encoding per edge:  hit_colors[2:0] =   
// 
//logic [0:15] [0:15] [2:0] hit_colors = 
//		  {48'o3333333333333333,     
//			48'o1333333333333332,    
//			48'o1133333333333322, 
//			48'o1113333333333222,
//			48'o1111333333332222,
//			48'o1111133333322222,
//			48'o1111113333222222,
//			48'o1111111332222222,
//			48'o1111111002222222,
//			48'o1111110000222222,
//			48'o1111100000022222,
//			48'o1111000000002222,
//			48'o1110000000000222,
//			48'o1100000000000022,
//			48'o1000000000000002,
//			48'o0000000000000000};
//			
//logic [0:15] [0:15] [2:0] hit_colors = 
//		  {48'o4433333333333344,     
//			48'o4443333333333444,    
//			48'o1444333333334442, 
//			48'o1144433333344422,
//			48'o1114443333444222,
//			48'o1111444334442222,
//			48'o1111144444422222,
//			48'o1111114444222222,
//			48'o1111114444222222,
//			48'o1111144444422222,
//			48'o1111444004442222,
//			48'o1114440000444222,
//			48'o1144400000044422,
//			48'o1444000000004442,
//			48'o4440000000000444,
//			48'o4400000000000044};


logic [0:3] [0:3] [3:0] hit_colors = 
			{16'h8442,
			 16'h8822,
			 16'h9933,
			 16'h9113};

 
 
// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		HitEdgeCode <= 3'h0;

	end

	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default  
		HitEdgeCode <= 3'h0;

		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket
		
			if (left_key)
				RGBout <= object_colors[1][offsetY][offsetX];
			else if (right_key)
				RGBout <= object_colors[1][offsetY][31 - offsetX];
			else if (up_key)
				RGBout <= object_colors[2][offsetY][offsetX];
			else
				RGBout <= object_colors[0][offsetY][offsetX];
			HitEdgeCode <= hit_colors[offsetY >> 3][offsetX >> 3];	//get hitting edge code from the colors table  
		
		end  	
	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule