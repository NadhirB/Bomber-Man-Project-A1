// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Feb 2025 
//(c) Technion IIT, Department of Electrical Engineering 2025 



module	WallsMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic col_blast_wall,
					input logic explosion,
					input logic game_on,
					input logic [3:0] layout_sel,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout    //rgb value from the bitmap
 ) ;
 

parameter int default_layout = 0;

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 


localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^5 = 32  everu object 
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 

localparam  int MAZE_NUMBER_OF__X_BITS = 5;  // 2^4 = 16 / /the maze of the objects 
localparam  int MAZE_NUMBER_OF__Y_BITS = 4;  // 2^3 = 8 

//-----

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;
localparam  int MAZE_WIDTH_X = 1 << MAZE_NUMBER_OF__X_BITS ;
localparam  int MAZE_HEIGHT_Y = 1 << MAZE_NUMBER_OF__Y_BITS ;


 logic [10:0] offsetX_LSB ;
 logic [10:0] offsetY_LSB ; 
 logic [10:0] offsetX_MSB ;
 logic [10:0] offsetY_MSB ;

 assign offsetX_LSB  = offsetX[(TILE_NUMBER_OF_X_BITS-1):0] ; // get lower bits 
 assign offsetY_LSB  = offsetY[(TILE_NUMBER_OF_Y_BITS-1):0] ; // get lower bits 
 assign offsetX_MSB  = offsetX[(TILE_NUMBER_OF_X_BITS + MAZE_NUMBER_OF__X_BITS -1 ):TILE_NUMBER_OF_X_BITS] ; // get higher bits 
 assign offsetY_MSB  = offsetY[(TILE_NUMBER_OF_Y_BITS + MAZE_NUMBER_OF__Y_BITS -1 ):TILE_NUMBER_OF_Y_BITS] ; // get higher bits 


 
// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 8 *16 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the understanding 



// This is a Test:

logic [1:0] MazeBitMapMask [0:12] [0:18];
logic MazeBitMapMask_exploding [0:12] [0:18];

logic [1:0] MazeDefaultBitMapMask [0:4] [0:12] [0:18] = 
		'{'{'{0, 3, 2, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0},
	  '{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1}, //col
	  '{0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 3, 1, 0, 0, 3, 3, 3, 1},
	  '{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0},
	  '{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1}, //col
	  '{0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 1},
	  '{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0},
	  '{0, 3, 0, 3, 0, 3, 3, 3, 0, 3, 0, 3, 0, 3, 3, 3, 1, 3, 1}, //col
	  '{0, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0},
	  '{2, 3, 2, 3, 0, 3, 3, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1}, //col
	  '{0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0}},
	  
		'{'{0, 0, 2, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0},
		'{0, 3, 0, 1, 0, 3, 0, 3, 1, 0, 0, 3, 0, 3, 1, 3, 0, 3, 1},
		'{0, 1, 0, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 3, 0, 1, 1},
		'{1, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 0, 0, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0},
		'{0, 3, 1, 0, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 0, 0, 3, 1},
		'{0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 3, 2, 0},
		'{0, 0, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 1, 0},
		'{0, 3, 0, 3, 3, 3, 0, 3, 0, 0, 0, 3, 1, 3, 3, 3, 1, 3, 1},
		'{0, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0},
		'{2, 3, 0, 0, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0}},
		
		'{'{0, 3, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1},
		'{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 1, 0, 1, 1, 1, 0, 0, 0, 1, 1, 2, 1, 0, 0, 3, 3, 0, 1},
		'{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0},
		'{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{1, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1},
		'{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 1},
		'{0, 3, 0, 3, 3, 3, 1, 3, 0, 3, 0, 3, 0, 3, 3, 3, 1, 3, 1},
		'{1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0},
		'{2, 3, 2, 3, 0, 3, 3, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1}},
		
		'{'{0, 0, 0, 0, 2, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 0, 0, 1},
		'{0, 3, 1, 3, 0, 0, 0, 3, 1, 3, 0, 3, 1, 3, 0, 0, 0, 3, 1},
		'{1, 0, 0, 1, 1, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 3, 1, 0},
		'{0, 3, 0, 0, 0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0},
		'{0, 3, 0, 3, 0, 3, 0, 0, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 1},
		'{0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0},
		'{0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 1, 0, 0, 0, 0, 0},
		'{0, 3, 0, 3, 3, 3, 1, 3, 0, 3, 0, 3, 0, 0, 3, 3, 1, 3, 1},
		'{0, 1, 0, 1, 1, 0, 1, 0, 1, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0},
		'{2, 3, 0, 3, 0, 3, 0, 0, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0}},
		
		
		'{'{0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 1, 0},
		'{0, 3, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 1, 3, 0, 0, 0, 3, 3, 0, 1},
		'{0, 3, 0, 3, 0, 3, 0, 0, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0},
		'{0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 0, 1, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1},
		'{0, 3, 0, 3, 0, 0, 0, 3, 0, 3, 0, 3, 1, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 1, 0, 0, 0, 0, 0},
		'{0, 3, 0, 3, 3, 3, 1, 3, 0, 3, 0, 3, 0, 3, 3, 3, 1, 3, 1},
		'{1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0},
		'{2, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 0, 3, 1},
		'{0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0}}
	  
	  };

logic MazeDefaultBitMapMask_exploding [0:12] [0:18] = 
	'{'{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}, //col
	  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}};
 
 


logic [0:2] [0:TILE_HEIGHT_Y-1] [0:TILE_WIDTH_X-1] [7:0] object_colors = {
	{{8'h6c,8'h6c,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h24},
	{8'h6c,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h24},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h24,8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'had,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h6c,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20},
	{8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20}},
	
	{{8'h6c,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h24},
	{8'h6c,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h24},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h00,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h20,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h20,8'h64,8'h64,8'h8c,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h6c,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h20,8'h20,8'h64,8'h00,8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h00,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'had,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h20,8'h64,8'h20,8'h20},
	{8'h8d,8'h20,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'had,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h20,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8c,8'h8c,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8c,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h00,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h20,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8c,8'h8c,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8c,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h20,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hb6,8'h20},
	{8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20}},
	
	{{8'h64,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h24},
	{8'h6c,8'h64,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h24,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h00,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h20,8'h64,8'h8c,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h8c,8'h20,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h20,8'h64,8'h20,8'h20,8'h20,8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h8d,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h20,8'h8d,8'h64,8'h84,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h8d,8'h64,8'h20,8'h00,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h8d,8'h8d,8'h20,8'h20,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h00,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h00,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'had,8'h64,8'h24,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h00,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h8d,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8c,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h20,8'h00,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8c,8'h8c,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h20,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h84,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h20,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h20,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8c,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20,8'h20,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h24,8'h20,8'h64,8'h20,8'h64,8'h64,8'h20,8'h64,8'h64,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h24,8'h20,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h20,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h00,8'h20,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h00,8'h20,8'h20,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20,8'h64,8'h64,8'h20,8'h20,8'h24,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h8d,8'h8d,8'h20,8'h20,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h6c,8'h20,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h64,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h20,8'h8d,8'h8d,8'h8d,8'h64,8'h20,8'h20,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h20,8'h64,8'h20,8'h8d,8'h8d,8'h20,8'h8d,8'h8d,8'h64,8'h20,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h20,8'h8d,8'h20,8'h8d,8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h20,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h24,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h20,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h8d,8'h8d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h20,8'h64,8'h64,8'h64,8'h64,8'h64,8'h20,8'h20},
	{8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hb6,8'h20},
	{8'h24,8'h24,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20}},
	
	};

 
//
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask[default_layout] ;  //  copy default tabel
		MazeBitMapMask_exploding <= MazeDefaultBitMapMask_exploding;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default
		if (!game_on) begin
			MazeBitMapMask <= MazeDefaultBitMapMask[layout_sel];
			end
		
		if (col_blast_wall) begin
			if (MazeBitMapMask[offsetY_MSB][offsetX_MSB] > 0 && MazeBitMapMask_exploding[offsetY_MSB][offsetX_MSB] != 1) begin
				MazeBitMapMask[offsetY_MSB][offsetX_MSB] <= MazeBitMapMask[offsetY_MSB][offsetX_MSB] - 1;
				MazeBitMapMask_exploding[offsetY_MSB][offsetX_MSB] <= 1;
			end
		end
		
		if (!explosion)
			MazeBitMapMask_exploding <= MazeDefaultBitMapMask_exploding;
		
		if (InsideRectangle == 1'b1 )	begin 
		   	case (MazeBitMapMask[offsetY_MSB][offsetX_MSB])
					 2'b00 : RGBout <= TRANSPARENT_ENCODING ;
					 2'b01 : RGBout <= object_colors[2][offsetY_LSB][offsetX_LSB];
					 2'b10 : RGBout <= object_colors[1][offsetY_LSB][offsetX_LSB];
					 2'b11 : RGBout <= object_colors[0][offsetY_LSB][offsetX_LSB];
				default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
				
			end
		

	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap 
endmodule

