// System-Verilog 'written by Alex Grinshpun May 2018
// New bitmap dudy February 2025
// (c) Technion IIT, Department of Electrical Engineering 2025 



module	playerBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic left_key,
					input logic right_key,
					input logic up_key,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
				   output   logic	[3:0] HitEdgeCode 
 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^5 = 32 


localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00;// RGB value in the bitmap representing a transparent pixel 

logic [0:2] [0:31] [0:31] [7:0] object_colors = {
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h46,8'h46,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h46,8'h46,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h65,8'h65,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h46,8'h46,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h46,8'h46,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h65,8'had,8'had,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'had,8'had,8'h65,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h65,8'had,8'had,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'had,8'had,8'h65,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h46,8'h46,8'hfa,8'hfa,8'hfa,8'hfa,8'h46,8'h46,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hd6,8'hd6,8'hfa,8'h46,8'h46,8'hfa,8'hfa,8'hfa,8'hfa,8'h46,8'h46,8'hfa,8'hd6,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hd6,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hc5,8'hc5,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hc5,8'hc5,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hfa,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'hfa,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hfa,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'hfa,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00},
	{8'h00,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h00},
	{8'h00,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h00},
	{8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00},
	{8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'h6d,8'h6d,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'hed,8'hed,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65},
	{8'h00,8'h65,8'h65,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'h65,8'h65},
	{8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h65,8'hc5,8'hc5,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hed,8'hc5,8'hc5,8'h65,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hfa,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'had,8'hfa,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'h65,8'h65,8'h65,8'had,8'had,8'had,8'h65,8'h65,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'hda,8'h65,8'h65,8'h65,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}}
	
	};


//////////--------------------------------------------------------------------------------------------------------------=



logic [0:7] [0:7] [3:0] hit_colors = 
			{32'hc4444446,
			 32'h8c444462,
			 32'h88c44622,
			 32'h888c6222,
			 32'h88893222,
			 32'h88911322,
			 32'h89111132,
			 32'h91111113};

 
 
// pipeline (ff) to get the pixel color from the array 	 

//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		HitEdgeCode <= 3'h0;

	end

	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default  
		HitEdgeCode <= 3'h0;

		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket
		
			//flip or cjange bitmap based on the direction the plyer is going in
			if (left_key)
				RGBout <= object_colors[1][offsetY][offsetX];
			else if (right_key)
				RGBout <= object_colors[1][offsetY][31 - offsetX];
			else if (up_key)
				RGBout <= object_colors[2][offsetY][offsetX];
			else
				RGBout <= object_colors[0][offsetY][offsetX];
			HitEdgeCode <= hit_colors[offsetY >> 2][offsetX >> 2];	//get hitting edge code from the colors table  
		
		end  	
	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 

always_comb 
begin
	
	drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap
	
end   

endmodule