
// This module holds all the bitmaps used for drawing the movment keys of the controls screen, both 1 and 2-player modes.



module	ControlsBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// o00set from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket

					output logic drawingRequest, //output that the pixel should be dispalyed 
					output logic [7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

 parameter int layout = 0;		// parameter to determind which key to display: 0 = 1-player, 1 = red player, 2 = blue player
 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 

localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^4 = 16  everu object 
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^4 = 16 

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;

 logic [10:0] offsetX_LSB  ;
 logic [10:0] offsetY_LSB  ; 
 logic [10:0] offsetX_MSB ;
 logic [10:0] offsetY_MSB  ;

 assign offsetX_LSB  = offsetX[(TILE_NUMBER_OF_X_BITS-1):0] ; // get lower bits 
 assign offsetY_LSB  = offsetY[(TILE_NUMBER_OF_Y_BITS-1):0] ; // get lower bits 
 assign offsetX_MSB  = offsetX[10:TILE_NUMBER_OF_X_BITS] ; // get higher bits 
 assign offsetY_MSB  = offsetY[10:TILE_NUMBER_OF_Y_BITS] ; // get higher bits 
 

 logic [0:10] [0:(TILE_HEIGHT_Y-1)][0:(TILE_WIDTH_X-1)] [7:0]  object_colors  = {
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'hda,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hba,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hda,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hb6,8'hff,8'hff,8'h71,8'h96,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h92,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hdf,8'hff,8'hff,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},


	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hda,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h96,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hba,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h96,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h96,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h92,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hba,8'hff,8'hff,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h96,8'h96,8'h96,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'hba,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hba,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h92,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h71,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hb6,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h91,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hdf,8'hff,8'hff,8'hb6,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hba,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hba,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hba,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'hda,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hba,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h96,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'hff,8'hff,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'hff,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}},
	
	
	{{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h96,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'h71,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'hff,8'hff,8'hff,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'hff,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h71,8'h71,8'hff,8'h71,8'hff,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'hff,8'hff,8'hff,8'h71,8'h71,8'hff,8'hff,8'h71,8'h71,8'h71,8'hff,8'hff,8'h71,8'hff,8'h71,8'hff,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h71,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}}
	
	
	
	
	
};
 
//
// pipeline (00) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
//		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		if (InsideRectangle == 1'b1 )	
			begin
			
			case (layout)
				0: begin
					case (offsetY_MSB)
					 0 : if (offsetX_MSB == 1) 
								RGBout <= object_colors[0][offsetY_LSB][offsetX_LSB] ;
							else
								RGBout <= TRANSPARENT_ENCODING ;
					 1 : if (offsetX_MSB == 0) 
								RGBout <= object_colors[1][offsetY_LSB][offsetX_LSB] ;
							else if (offsetX_MSB == 1)
								RGBout <= object_colors[2][offsetY_LSB][offsetX_LSB] ; 
							else if (offsetX_MSB == 2)
								RGBout <= object_colors[3][offsetY_LSB][offsetX_LSB] ;
							else
								RGBout <= TRANSPARENT_ENCODING ;
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
				
				end
				
				1: begin
					case (offsetY_MSB)
					 0 : if (offsetX_MSB == 1) 
								RGBout <= object_colors[5][offsetY_LSB][offsetX_LSB] ;
							else
								RGBout <= TRANSPARENT_ENCODING ;
					 1 : if (offsetX_MSB == 0) 
								RGBout <= object_colors[4][offsetY_LSB][offsetX_LSB] ;
							else if (offsetX_MSB == 1)
								RGBout <= object_colors[6][offsetY_LSB][offsetX_LSB] ; 
							else if (offsetX_MSB == 2)
								RGBout <= object_colors[7][offsetY_LSB][offsetX_LSB] ;
							else
								RGBout <= TRANSPARENT_ENCODING ;
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
				
				end
				
				
				2: begin
					case (offsetY_MSB)
					 0 : if (offsetX_MSB == 1) 
								RGBout <= object_colors[0][offsetY_LSB][offsetX_LSB] ;
							else
								RGBout <= TRANSPARENT_ENCODING ;
					 1 : if (offsetX_MSB == 0) 
								RGBout <= object_colors[9][offsetY_LSB][offsetX_LSB] ;
							else if (offsetX_MSB == 1)
								RGBout <= object_colors[8][offsetY_LSB][offsetX_LSB] ; 
							else if (offsetX_MSB == 2)
								RGBout <= object_colors[10][offsetY_LSB][offsetX_LSB] ;
							else
								RGBout <= TRANSPARENT_ENCODING ;
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
				
				end
				
				
				default: RGBout <= TRANSPARENT_ENCODING;
			
			
			endcase
			end 
		

	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

