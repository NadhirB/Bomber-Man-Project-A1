// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Feb 2025 
//(c) Technion IIT, Department of Electrical Engineering 2025 



module	blueblastMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket
					input logic [2:0] blast_num,
					input logic blast,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 


localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^5 = 32  everu object 
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 

localparam  int MAZE_NUMBER_OF__X_BITS = 4;  // 2^4 = 16 / /the maze of the objects 
localparam  int MAZE_NUMBER_OF__Y_BITS = 3;  // 2^3 = 8 

//-----

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;
localparam  int MAZE_WIDTH_X = 1 << MAZE_NUMBER_OF__X_BITS ;
localparam  int MAZE_HEIGHT_Y = 1 << MAZE_NUMBER_OF__Y_BITS ;


 logic [10:0] offsetX_LSB  ;
 logic [10:0] offsetY_LSB  ; 
 logic [10:0] offsetX_MSB ;
 logic [10:0] offsetY_MSB  ;
 logic [2:0] blast_num_D;

 assign offsetX_LSB  = offsetX[(TILE_NUMBER_OF_X_BITS-1):0] ; // get lower bits 
 assign offsetY_LSB  = offsetY[(TILE_NUMBER_OF_Y_BITS-1):0] ; // get lower bits 
 assign offsetX_MSB  = offsetX[(TILE_NUMBER_OF_X_BITS + MAZE_NUMBER_OF__X_BITS -1 ):TILE_NUMBER_OF_X_BITS] ; // get higher bits 
 assign offsetY_MSB  = offsetY[(TILE_NUMBER_OF_Y_BITS + MAZE_NUMBER_OF__Y_BITS -1 ):TILE_NUMBER_OF_Y_BITS] ; // get higher bits 
 

 
// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 8 *16 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the understanding 



// This is a Test:

logic [1:0] MazeBitMapMask [0:2] [0:4] [0:4];

logic [1:0] MazeDefaultBitMapMask [0:2] [0:4] [0:4] = '{
	'{'{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b1, 1'b1, 1'b1, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0}},
	  
	'{'{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b1, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0}},
	  
	'{'{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b1, 1'b1, 1'b1, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
	  '{1'b0, 1'b0, 1'b0, 1'b0, 1'b0}}};
 

logic [0:TILE_HEIGHT_Y-1] [0:TILE_WIDTH_X-1] [7:0] object_colors = {
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h25,8'h25,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h26,8'hFF,8'hFF,8'h05,8'hFF,8'h05,8'h06,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h2f,8'h2f,8'h26,8'hFF,8'h05,8'hFF,8'h06,8'hFF,8'h2f,8'hFF,8'hFF,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'hFF,8'hFF,8'hFF,8'h2f,8'h1b,8'h27,8'h2f,8'h25,8'h25,8'h05,8'h05,8'h2f,8'h1b,8'h25,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h01,8'h26,8'h05,8'h26,8'hFF,8'hFF,8'h1b,8'h7f,8'h1b,8'h1b,8'h05,8'h2f,8'h2f,8'h1b,8'hdf,8'h05,8'hFF,8'hFF,8'h26,8'h05,8'h26,8'h25,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h2e,8'h05,8'h25,8'h05,8'h05,8'h2d,8'hdf,8'h3f,8'h1b,8'h2f,8'h2f,8'h2f,8'h1b,8'hdf,8'h25,8'h05,8'h05,8'h05,8'h05,8'h26,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h26,8'h25,8'h25,8'h05,8'h2f,8'h1b,8'hbf,8'h3f,8'hdf,8'h1b,8'h2f,8'h3f,8'hdf,8'h1b,8'h2f,8'h2f,8'h05,8'h05,8'h25,8'h26,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'h2f,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h05,8'h25,8'h25,8'h2f,8'h26,8'h1b,8'hdf,8'hbf,8'h1b,8'hbf,8'h1b,8'h1b,8'h2f,8'h25,8'h05,8'h2e,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'h3f,8'h2f,8'h33,8'h05,8'h05,8'h05,8'h2f,8'h25,8'h05,8'h2f,8'h1b,8'hdf,8'hdf,8'hdf,8'hdf,8'h27,8'h3f,8'h1b,8'h25,8'h25,8'h2f,8'h2f,8'h05,8'hFF,8'h2f,8'h2f,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h1b,8'h2f,8'h1b,8'h25,8'h1f,8'h25,8'h25,8'hbf,8'h2f,8'h3f,8'h1b,8'h3f,8'h33,8'h1b,8'hdf,8'h25,8'h2f,8'h2f,8'h1b,8'h1b,8'hbf,8'h2f,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'h2f,8'h1b,8'h1b,8'hdf,8'hdf,8'h1f,8'h1b,8'hdf,8'h1b,8'h33,8'h33,8'h1b,8'h33,8'h3f,8'hdf,8'h3f,8'hdf,8'h2f,8'h25,8'hdf,8'hdf,8'h3f,8'h25,8'h2f,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'h05,8'h05,8'h05,8'h2f,8'h1b,8'h9f,8'h1f,8'h1f,8'h1f,8'hdf,8'h3f,8'hbf,8'h3f,8'h3f,8'h3f,8'h3f,8'h2f,8'h2f,8'hdf,8'h3f,8'h1b,8'h3f,8'h2f,8'h2f,8'hFF,8'h05,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h05,8'h2f,8'h33,8'h3f,8'h2f,8'h1b,8'h9f,8'h1b,8'hdf,8'hdf,8'hdf,8'hdf,8'hbf,8'h1b,8'h3f,8'hdf,8'hdf,8'hdf,8'h2f,8'h2f,8'h05,8'h05,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'h05,8'h26,8'h05,8'h05,8'h05,8'h2f,8'h2f,8'h1b,8'h1f,8'hdf,8'h3f,8'h1b,8'h3f,8'hdf,8'hdf,8'hdf,8'h3f,8'h3f,8'h1b,8'h37,8'h7f,8'hdf,8'h3f,8'h2f,8'h25,8'h2f,8'h05,8'h05,8'h26,8'h25,8'hFF},
	{8'hFF,8'h25,8'h26,8'h05,8'h05,8'h2f,8'h25,8'h2f,8'h3b,8'hdf,8'h3f,8'h37,8'h1b,8'h3f,8'h3f,8'hdf,8'hdf,8'hdf,8'h3f,8'h1b,8'hbf,8'hdf,8'h1b,8'h1b,8'h2f,8'h2f,8'h05,8'h05,8'h05,8'h26,8'h25,8'hFF},
	{8'hFF,8'hFF,8'h01,8'hFF,8'h05,8'h05,8'h2f,8'h2f,8'hdf,8'hdf,8'hdf,8'h1f,8'h3b,8'hbf,8'hdf,8'hdf,8'h7f,8'hdf,8'h3f,8'hbf,8'h1b,8'h2f,8'h3f,8'h33,8'h2f,8'h05,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'h01,8'hFF,8'h2f,8'h2f,8'h3f,8'h3f,8'h3f,8'hdf,8'h2f,8'h2f,8'h3f,8'h3f,8'h3f,8'h3f,8'h9f,8'h3f,8'hdf,8'h3b,8'h3f,8'h3f,8'h7f,8'h1b,8'h17,8'h05,8'h05,8'h01,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'h2f,8'h25,8'h1f,8'hdf,8'hdf,8'h25,8'h2f,8'h9f,8'h3f,8'hdf,8'h3f,8'h33,8'h1b,8'h33,8'h2f,8'h1b,8'hdf,8'h1b,8'h1f,8'hdf,8'hdf,8'h1b,8'h1b,8'h2f,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h2f,8'hdf,8'h1b,8'h2e,8'h2f,8'h2f,8'h25,8'hbf,8'h3b,8'h33,8'h3f,8'h1b,8'h3f,8'h2f,8'hdf,8'h05,8'h25,8'h1b,8'h2f,8'h3f,8'h2f,8'h1b,8'h27,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'h26,8'h2f,8'hFF,8'h05,8'h2f,8'h2f,8'h25,8'h05,8'h1b,8'h3f,8'h2f,8'hdf,8'hbf,8'hdf,8'hbf,8'h1b,8'h2f,8'h05,8'h06,8'h2f,8'h05,8'h05,8'h05,8'h2f,8'h2f,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h25,8'h05,8'h26,8'h2f,8'h1b,8'h1b,8'hdf,8'h1b,8'hbf,8'hdf,8'h1f,8'h2f,8'h2f,8'h25,8'h25,8'h05,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h06,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h2e,8'h2e,8'h25,8'h05,8'h2f,8'h2f,8'h37,8'hdf,8'h3f,8'h2f,8'h1b,8'hdf,8'h3f,8'hdf,8'h1b,8'h2f,8'h25,8'h05,8'h05,8'h26,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h05,8'h25,8'h05,8'h05,8'h25,8'hbf,8'h1b,8'h2f,8'h33,8'h2f,8'h33,8'h3f,8'hdf,8'h27,8'h05,8'h05,8'h05,8'h05,8'h26,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h01,8'h2e,8'h25,8'h25,8'hFF,8'hFF,8'h05,8'h9f,8'h1b,8'h2f,8'h2f,8'h05,8'h1b,8'h1b,8'h3f,8'h1b,8'hFF,8'hFF,8'h25,8'h25,8'h05,8'h25,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'h25,8'h1b,8'h2f,8'h05,8'h05,8'h2e,8'h25,8'h2f,8'h2f,8'h3f,8'h06,8'hFF,8'hFF,8'hFF,8'h25,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'hFF,8'hFF,8'h2f,8'hFF,8'h05,8'hFF,8'h05,8'hFF,8'h2f,8'h2f,8'h2f,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h06,8'hFF,8'h05,8'hFF,8'hFF,8'h26,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h25,8'h26,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h05,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}};

 
//
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
		blast_num_D <= 0;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		
		if (!blast)
			blast_num_D <= blast_num;
			
		if (InsideRectangle == 1'b1 )	
			begin 
		   	case (MazeBitMapMask[blast_num_D][offsetY_MSB][offsetX_MSB])
					 1'b0 : RGBout <= TRANSPARENT_ENCODING ;
					 1'b1 : RGBout <= object_colors[offsetY_LSB][offsetX_LSB];  
				default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
			end 

	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

