

module	DoorIdolBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic select,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout    //rgb value from the bitmap
 ) ;
 


localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^5 = 32  everu object 
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 


//-----

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h01 ;// RGB value in the bitmap representing a transparent pixel 

logic [0:1] [0:TILE_HEIGHT_Y-1] [0:TILE_WIDTH_X-1] [7:0] object_colors = {
	{{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'hdf,8'hdf,8'hdf,8'hdf,8'h72,8'h6d,8'h6d,8'h72,8'h6d,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h6d,8'h72,8'h6d,8'h6d,8'h72,8'hdf,8'hdf,8'hdf,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h64,8'h64,8'h6d,8'h6d,8'h72,8'h6d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h6d,8'h72,8'h6d,8'h6d,8'h64,8'h64,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h64,8'h64,8'h6d,8'h6d,8'h72,8'h6d,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h6d,8'h72,8'h6d,8'h6d,8'h64,8'h64,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h6d,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'hb1,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'hb1,8'h64,8'h6d,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'hb1,8'hb1,8'hb1,8'h64,8'h6d,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h6d,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h91,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'h91,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h6d,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'hb1,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h6d,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'hb1,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'h64,8'h64,8'hb1,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'hb1,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'hb1,8'h64,8'h64,8'hb1,8'h6d,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'h6d,8'h6d,8'h64,8'h6d,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'h6d,8'h6d,8'h6d,8'h64,8'h6d,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'h72,8'hdf,8'hdf,8'hdf,8'hdf,8'h72,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'hb1,8'h72,8'hdf,8'hdf,8'hdf,8'hdf,8'h72,8'hb1,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'h72,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'hb1,8'hb1,8'h64,8'h64,8'h6d,8'h72,8'hdf,8'hdf,8'hdf,8'hdf,8'h72,8'h6d,8'h64,8'h64,8'hb1,8'hb1,8'hb1,8'hb1,8'h64,8'hb1,8'h64,8'h64,8'h72,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h6d,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h64,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h6d,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'h64,8'hdf,8'h6d},
	{8'h6d,8'hdf,8'hdf,8'hdf,8'hdf,8'h72,8'hdf,8'hdf,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'hdf,8'hdf,8'h72,8'hdf,8'hdf,8'hdf,8'hdf,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d}},
	
	{{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h00,8'h20,8'h20,8'h20,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h20,8'h20,8'h20,8'h00,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h00,8'h20,8'h20,8'h20,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h20,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h84,8'hf0,8'hf0,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h84,8'hf0,8'hf0,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfd,8'hfd,8'hf0,8'hf0,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'hf0,8'hf0,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfd,8'hfd,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'hf0,8'hfd,8'hf0,8'h20,8'h20,8'h84,8'h84,8'hf0,8'hf0,8'hf0,8'hf0,8'h84,8'h84,8'h20,8'h20,8'hf0,8'hfd,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'h84,8'hf0,8'h20,8'h20,8'h20,8'h20,8'h84,8'hf0,8'hf4,8'hf4,8'hf0,8'h84,8'h20,8'h20,8'h20,8'h20,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'h84,8'hf0,8'h84,8'h84,8'h20,8'h20,8'hf0,8'hf4,8'hff,8'hff,8'hf4,8'hf0,8'h20,8'h20,8'h84,8'h84,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'h84,8'hf0,8'hfd,8'hf0,8'h84,8'h84,8'h20,8'hf4,8'hfd,8'hff,8'hff,8'hfd,8'hf4,8'h20,8'h84,8'h84,8'hf0,8'hfd,8'h84,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'hf0,8'hf4,8'hff,8'hff,8'hf0,8'hf0,8'hf0,8'hfd,8'hfd,8'hff,8'hff,8'hfd,8'hfd,8'hf0,8'hf0,8'hf0,8'hff,8'hff,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h00,8'h84,8'hff,8'h84,8'hf4,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hf0,8'hfd,8'hfd,8'hff,8'hff,8'hfd,8'hfd,8'hf0,8'hff,8'hff,8'hff,8'hff,8'hf4,8'h84,8'hff,8'h84,8'h00,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h00,8'h84,8'hff,8'h84,8'hf4,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'h84,8'h20,8'h84,8'h84,8'h20,8'h84,8'hf0,8'hfd,8'hfd,8'hfd,8'hfd,8'hf4,8'h84,8'hff,8'h84,8'h00,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h00,8'h84,8'hfd,8'h84,8'hf4,8'hf4,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'hf0,8'h20,8'h84,8'h84,8'h20,8'hf0,8'hf0,8'hfd,8'hfd,8'hfd,8'hfd,8'hf4,8'h84,8'hfd,8'h84,8'h00,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h00,8'h84,8'hf0,8'hf0,8'hf4,8'hf4,8'hf0,8'h84,8'h84,8'hf0,8'h20,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'h20,8'hf0,8'h84,8'h84,8'hf0,8'hf4,8'hf0,8'hf0,8'h84,8'h00,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h00,8'h20,8'h84,8'hf0,8'hf4,8'hf0,8'h84,8'h84,8'h84,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h84,8'h84,8'h84,8'hf4,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h00,8'h20,8'h20,8'h84,8'hf0,8'h84,8'h84,8'h84,8'h20,8'h20,8'hf0,8'hf0,8'h20,8'hf0,8'hf0,8'h20,8'hf0,8'hf0,8'h20,8'h20,8'h84,8'h84,8'hf0,8'h84,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h84,8'h84,8'h84,8'h20,8'h84,8'h20,8'h84,8'hf0,8'h20,8'hfd,8'hfd,8'h20,8'hf0,8'h84,8'h20,8'h84,8'h20,8'h84,8'h84,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h20,8'h84,8'hf0,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hf0,8'h20,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'h20,8'hf0,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'hf0,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h20,8'hf0,8'h20,8'h84,8'h20,8'h84,8'hf0,8'h20,8'hfd,8'hfd,8'h20,8'hf0,8'h84,8'h20,8'h84,8'h20,8'hf0,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'h20,8'hfc,8'hfc,8'h84,8'h20,8'hf0,8'hf0,8'h20,8'hf0,8'hf0,8'h20,8'hf0,8'hf0,8'h20,8'h84,8'hfc,8'hfc,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h20,8'hf4,8'hf4,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hf4,8'hf4,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h84,8'h20,8'hf4,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hf4,8'h20,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'h84,8'h20,8'h84,8'h84,8'hf0,8'hf0,8'hfd,8'hfd,8'hfd,8'hfd,8'hf0,8'hf0,8'h84,8'h84,8'h20,8'h84,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'hf0,8'hf0,8'hf0,8'hfc,8'hfc,8'hff,8'hff,8'hf0,8'hf0,8'hf0,8'hf0,8'hff,8'hff,8'hfc,8'hfc,8'hf0,8'hf0,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h84,8'hf0,8'hf0,8'hfc,8'hfc,8'hfc,8'hfc,8'hff,8'hf0,8'hf0,8'hff,8'hfc,8'hfc,8'hfc,8'hfc,8'hf0,8'hf0,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h20,8'hf0,8'hf0,8'hf0,8'hf0,8'h84,8'h84,8'h84,8'h84,8'hf0,8'hf0,8'hf0,8'hf0,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h20,8'h20,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h84,8'h20,8'h20,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01}}
	
	};

 
//
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default
		
		
		if (InsideRectangle == 1'b1 )	begin 
		   RGBout <= object_colors[select][offsetY][offsetX];
			end
		

	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap 
endmodule

